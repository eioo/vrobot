module vrobot

struct Color {
pub:
  r int
  g int
  b int
}

struct Size {
pub:
  width int
  height int
}

struct Point {
pub:
  x int
  y int
}
