module vrobot
 
#flag -lgdi32
#include "windows.h"
