module vrobot
 
import math
import time

#flag -lgdi32
#include "windows.h"
