module vrobot

struct Color {
pub:
  r int
  g int
  b int
}

struct Point {
pub:
  x int
  y int
}
